/*
 * Experiments with loop constructs in SV. Refer Section 12 of 2012 LRM
 * 
 */

module loops();

   int sampleA_unpkd [10] = '{0,1,2,3,4,5,6,7,8,9};
   int sampleB[4];

   
   
endmodule : loops

